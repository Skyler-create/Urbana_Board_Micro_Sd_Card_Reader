module color_mapper(


);

endmodule